magic
tech sky130A
timestamp 1725643987
<< nwell >>
rect -168 121 53 352
rect 180 121 401 352
rect 528 132 735 348
<< nmos >>
rect -24 -13 -9 87
rect 324 -13 339 87
rect 662 12 677 72
<< pmos >>
rect -24 139 -9 334
rect 324 139 339 334
rect 662 150 677 330
<< ndiff >>
rect -56 58 -24 87
rect -56 7 -52 58
rect -35 7 -24 58
rect -56 -13 -24 7
rect -9 62 23 87
rect -9 11 2 62
rect 19 11 23 62
rect -9 -13 23 11
rect 292 58 324 87
rect 292 7 296 58
rect 313 7 324 58
rect 292 -13 324 7
rect 339 62 371 87
rect 339 11 350 62
rect 367 11 371 62
rect 625 60 662 72
rect 625 24 633 60
rect 653 24 662 60
rect 625 12 662 24
rect 677 59 712 72
rect 677 23 688 59
rect 708 23 712 59
rect 677 12 712 23
rect 339 -13 371 11
<< pdiff >>
rect -63 281 -24 334
rect -63 219 -55 281
rect -38 219 -24 281
rect -63 139 -24 219
rect -9 250 30 334
rect -9 188 3 250
rect 20 188 30 250
rect -9 139 30 188
rect 285 281 324 334
rect 285 219 293 281
rect 310 219 324 281
rect 285 139 324 219
rect 339 250 378 334
rect 339 188 351 250
rect 368 188 378 250
rect 339 139 378 188
rect 622 294 662 330
rect 622 180 628 294
rect 651 180 662 294
rect 622 150 662 180
rect 677 294 717 330
rect 677 180 686 294
rect 709 180 717 294
rect 677 150 717 180
<< ndiffc >>
rect -52 7 -35 58
rect 2 11 19 62
rect 296 7 313 58
rect 350 11 367 62
rect 633 24 653 60
rect 688 23 708 59
<< pdiffc >>
rect -55 219 -38 281
rect 3 188 20 250
rect 293 219 310 281
rect 351 188 368 250
rect 628 180 651 294
rect 686 180 709 294
<< psubdiff >>
rect -117 57 -56 87
rect -117 7 -108 57
rect -83 7 -56 57
rect -117 -13 -56 7
rect 231 51 292 87
rect 231 1 240 51
rect 265 1 292 51
rect 231 -13 292 1
rect 554 60 625 72
rect 554 22 575 60
rect 598 22 625 60
rect 554 12 625 22
<< nsubdiff >>
rect -150 304 -63 334
rect -150 217 -141 304
rect -112 217 -63 304
rect -150 139 -63 217
rect 198 318 285 334
rect 198 229 206 318
rect 231 229 285 318
rect 198 139 285 229
rect 546 294 622 330
rect 546 179 562 294
rect 601 179 622 294
rect 546 150 622 179
<< psubdiffcont >>
rect -108 7 -83 57
rect 240 1 265 51
rect 575 22 598 60
<< nsubdiffcont >>
rect -141 217 -112 304
rect 206 229 231 318
rect 562 179 601 294
<< poly >>
rect -24 334 -9 347
rect 324 334 339 347
rect 662 330 677 347
rect -24 87 -9 139
rect 324 87 339 139
rect 461 128 499 134
rect 662 128 677 150
rect 461 124 677 128
rect 461 106 470 124
rect 487 106 677 124
rect 461 102 677 106
rect 461 97 505 102
rect 662 72 677 102
rect -24 -67 -9 -13
rect 324 -67 339 -13
rect 662 -25 677 12
<< polycont >>
rect 470 106 487 124
<< locali >>
rect 285 451 315 452
rect -169 447 694 451
rect -169 424 -145 447
rect -113 444 694 447
rect -113 424 79 444
rect -169 421 79 424
rect 111 443 694 444
rect 111 421 306 443
rect -169 420 306 421
rect 338 420 580 443
rect 612 420 694 443
rect -169 408 694 420
rect -150 304 -101 408
rect -150 217 -141 304
rect -112 217 -101 304
rect -150 200 -101 217
rect -63 281 -33 408
rect -63 219 -55 281
rect -38 219 -33 281
rect 198 318 240 408
rect -63 200 -33 219
rect -2 250 25 267
rect -2 188 3 250
rect 20 188 25 250
rect 198 229 206 318
rect 231 229 240 318
rect 198 207 240 229
rect 285 281 315 408
rect 562 306 607 408
rect 285 219 293 281
rect 310 219 315 281
rect 550 294 658 306
rect 285 207 315 219
rect 346 250 373 267
rect -2 172 25 188
rect 346 188 351 250
rect 368 188 373 250
rect 346 172 373 188
rect 550 179 562 294
rect 601 180 628 294
rect 651 180 658 294
rect 601 179 658 180
rect -2 155 490 172
rect 550 163 658 179
rect 681 294 714 306
rect 681 180 686 294
rect 709 180 714 294
rect 681 163 714 180
rect -117 57 -76 78
rect -117 7 -108 57
rect -83 7 -76 57
rect -117 -4 -76 7
rect -56 58 -31 78
rect -56 7 -52 58
rect -35 7 -31 58
rect -116 -97 -78 -4
rect -56 -30 -31 7
rect -2 62 23 155
rect 462 134 490 155
rect 462 124 499 134
rect -2 11 2 62
rect 19 11 23 62
rect -2 -4 23 11
rect 181 94 371 112
rect 462 106 470 124
rect 487 106 499 124
rect 462 102 499 106
rect 181 -30 212 94
rect 292 60 317 77
rect 231 58 317 60
rect 231 51 296 58
rect 231 1 240 51
rect 265 7 296 51
rect 313 7 317 58
rect 265 1 317 7
rect 231 -4 317 1
rect 346 62 371 94
rect 346 11 350 62
rect 367 11 371 62
rect 567 60 656 68
rect 686 67 707 163
rect 567 22 575 60
rect 598 24 633 60
rect 653 24 656 60
rect 598 22 656 24
rect 567 15 656 22
rect 683 59 710 67
rect 683 23 688 59
rect 708 23 710 59
rect 683 15 710 23
rect 231 -7 269 -4
rect -56 -47 212 -30
rect 237 -97 268 -7
rect 346 -9 371 11
rect 573 -97 615 15
rect -182 -103 681 -97
rect -182 -108 101 -103
rect -182 -133 -156 -108
rect -115 -128 101 -108
rect 142 -106 681 -103
rect 142 -128 341 -106
rect -115 -131 341 -128
rect 382 -107 681 -106
rect 382 -131 589 -107
rect -115 -132 589 -131
rect 630 -132 681 -107
rect -115 -133 681 -132
rect -182 -145 681 -133
<< viali >>
rect -145 424 -113 447
rect 79 421 111 444
rect 306 420 338 443
rect 580 420 612 443
rect -156 -133 -115 -108
rect 101 -128 142 -103
rect 341 -131 382 -106
rect 589 -132 630 -107
<< metal1 >>
rect -172 447 698 453
rect -172 424 -145 447
rect -113 444 698 447
rect -113 424 79 444
rect -172 421 79 424
rect 111 443 698 444
rect 111 421 306 443
rect -172 420 306 421
rect 338 420 580 443
rect 612 420 698 443
rect -172 399 698 420
rect -189 -103 681 -91
rect -189 -108 101 -103
rect -189 -133 -156 -108
rect -115 -128 101 -108
rect 142 -106 681 -103
rect 142 -128 341 -106
rect -115 -131 341 -128
rect 382 -107 681 -106
rect 382 -131 589 -107
rect -115 -132 589 -131
rect 630 -132 681 -107
rect -115 -133 681 -132
rect -189 -145 681 -133
<< labels >>
flabel poly -16 -49 -16 -49 0 FreeSans 40 0 0 0 c
port 0 nsew
flabel poly 331 -53 331 -53 0 FreeSans 40 0 0 0 d
port 1 nsew
flabel locali 696 111 696 111 0 FreeSans 40 0 0 0 out
port 2 nsew
flabel metal1 243 431 243 431 0 FreeSans 40 0 0 0 vdd
port 3 nsew
flabel metal1 266 -126 266 -126 0 FreeSans 40 0 0 0 vss
port 5 nsew
<< end >>
