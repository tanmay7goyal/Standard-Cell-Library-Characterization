magic
tech sky130A
timestamp 1726334538
<< nwell >>
rect 2710 345 2827 346
rect -892 118 -678 312
rect -487 118 -273 312
rect -85 106 124 324
rect 263 118 477 312
rect 611 118 825 312
rect 1061 117 1294 335
rect 1564 106 1773 324
rect 1912 118 2126 312
rect 2260 118 2474 312
rect 2710 127 2943 345
rect 3162 118 3376 312
<< nmos >>
rect 20 1 35 61
rect -759 -97 -744 -55
rect -354 -97 -339 -55
rect 744 -45 759 -3
rect 396 -97 411 -55
rect 1190 -55 1205 5
rect 1669 -62 1684 -2
rect 2393 -45 2408 -3
rect 2045 -97 2060 -55
rect 2839 -55 2854 5
rect 3295 -97 3310 -55
<< pmos >>
rect -759 150 -744 285
rect -354 150 -339 285
rect 20 126 35 306
rect 396 150 411 285
rect 744 150 759 285
rect 1190 137 1205 317
rect 1669 126 1684 306
rect 2045 150 2060 285
rect 2393 150 2408 285
rect 2839 147 2854 327
rect 3295 150 3310 285
<< ndiff >>
rect -10 41 20 61
rect -10 11 -6 41
rect 14 11 20 41
rect -10 1 20 11
rect 35 41 70 61
rect 35 11 45 41
rect 65 11 70 41
rect 35 1 70 11
rect -802 -62 -759 -55
rect -802 -87 -794 -62
rect -776 -87 -759 -62
rect -802 -97 -759 -87
rect -744 -62 -704 -55
rect -744 -87 -731 -62
rect -713 -87 -704 -62
rect -744 -97 -704 -87
rect -397 -62 -354 -55
rect -397 -87 -389 -62
rect -371 -87 -354 -62
rect -397 -97 -354 -87
rect -339 -62 -299 -55
rect 701 -10 744 -3
rect 701 -35 709 -10
rect 727 -35 744 -10
rect 701 -45 744 -35
rect 759 -10 832 -3
rect 759 -35 805 -10
rect 823 -35 832 -10
rect 759 -45 832 -35
rect 1160 -15 1190 5
rect -339 -87 -326 -62
rect -308 -87 -299 -62
rect -339 -97 -299 -87
rect 353 -62 396 -55
rect 353 -87 361 -62
rect 379 -87 396 -62
rect 353 -97 396 -87
rect 411 -62 451 -55
rect 411 -87 424 -62
rect 442 -87 451 -62
rect 1160 -45 1164 -15
rect 1184 -45 1190 -15
rect 1160 -55 1190 -45
rect 1205 -15 1240 5
rect 1205 -45 1215 -15
rect 1235 -45 1240 -15
rect 1639 -22 1669 -2
rect 1205 -55 1240 -45
rect 1639 -52 1643 -22
rect 1663 -52 1669 -22
rect 1639 -62 1669 -52
rect 1684 -22 1719 -2
rect 1684 -52 1694 -22
rect 1714 -52 1719 -22
rect 1684 -62 1719 -52
rect 2350 -10 2393 -3
rect 2350 -35 2358 -10
rect 2376 -35 2393 -10
rect 2350 -45 2393 -35
rect 2408 -10 2481 -3
rect 2408 -35 2454 -10
rect 2472 -35 2481 -10
rect 2408 -45 2481 -35
rect 2809 -15 2839 5
rect 2002 -62 2045 -55
rect 411 -97 451 -87
rect 2002 -87 2010 -62
rect 2028 -87 2045 -62
rect 2002 -97 2045 -87
rect 2060 -62 2100 -55
rect 2060 -87 2073 -62
rect 2091 -87 2100 -62
rect 2809 -45 2813 -15
rect 2833 -45 2839 -15
rect 2809 -55 2839 -45
rect 2854 -15 2889 5
rect 2854 -45 2864 -15
rect 2884 -45 2889 -15
rect 2854 -55 2889 -45
rect 3252 -62 3295 -55
rect 2060 -97 2100 -87
rect 3252 -87 3260 -62
rect 3278 -87 3295 -62
rect 3252 -97 3295 -87
rect 3310 -62 3350 -55
rect 3310 -87 3323 -62
rect 3341 -87 3350 -62
rect 3310 -97 3350 -87
<< pdiff >>
rect -832 273 -759 285
rect -832 248 -823 273
rect -805 248 -759 273
rect -832 150 -759 248
rect -744 185 -704 285
rect -744 160 -731 185
rect -713 160 -704 185
rect -744 150 -704 160
rect -427 273 -354 285
rect -427 248 -418 273
rect -400 248 -354 273
rect -427 150 -354 248
rect -339 185 -299 285
rect -339 160 -326 185
rect -308 160 -299 185
rect -339 150 -299 160
rect -10 166 20 306
rect -10 136 -6 166
rect 14 136 20 166
rect -10 126 20 136
rect 35 166 70 306
rect 35 136 45 166
rect 65 136 70 166
rect 323 273 396 285
rect 323 248 332 273
rect 350 248 396 273
rect 323 150 396 248
rect 411 185 451 285
rect 411 160 424 185
rect 442 160 451 185
rect 411 150 451 160
rect 671 273 744 285
rect 671 248 680 273
rect 698 248 744 273
rect 671 150 744 248
rect 759 185 799 285
rect 759 160 772 185
rect 790 160 799 185
rect 759 150 799 160
rect 35 126 70 136
rect 1160 177 1190 317
rect 1160 147 1164 177
rect 1184 147 1190 177
rect 1160 137 1190 147
rect 1205 177 1240 317
rect 1205 147 1215 177
rect 1235 147 1240 177
rect 1205 137 1240 147
rect 1639 166 1669 306
rect 1639 136 1643 166
rect 1663 136 1669 166
rect 1639 126 1669 136
rect 1684 166 1719 306
rect 1684 136 1694 166
rect 1714 136 1719 166
rect 1972 273 2045 285
rect 1972 248 1981 273
rect 1999 248 2045 273
rect 1972 150 2045 248
rect 2060 185 2100 285
rect 2060 160 2073 185
rect 2091 160 2100 185
rect 2060 150 2100 160
rect 2320 273 2393 285
rect 2320 248 2329 273
rect 2347 248 2393 273
rect 2320 150 2393 248
rect 2408 185 2448 285
rect 2408 160 2421 185
rect 2439 160 2448 185
rect 2408 150 2448 160
rect 1684 126 1719 136
rect 2809 187 2839 327
rect 2809 157 2813 187
rect 2833 157 2839 187
rect 2809 147 2839 157
rect 2854 187 2889 327
rect 2854 157 2864 187
rect 2884 157 2889 187
rect 2854 147 2889 157
rect 3222 273 3295 285
rect 3222 248 3231 273
rect 3249 248 3295 273
rect 3222 150 3295 248
rect 3310 185 3350 285
rect 3310 160 3323 185
rect 3341 160 3350 185
rect 3310 150 3350 160
<< ndiffc >>
rect -6 11 14 41
rect 45 11 65 41
rect -794 -87 -776 -62
rect -731 -87 -713 -62
rect -389 -87 -371 -62
rect 709 -35 727 -10
rect 805 -35 823 -10
rect -326 -87 -308 -62
rect 361 -87 379 -62
rect 424 -87 442 -62
rect 1164 -45 1184 -15
rect 1215 -45 1235 -15
rect 1643 -52 1663 -22
rect 1694 -52 1714 -22
rect 2358 -35 2376 -10
rect 2454 -35 2472 -10
rect 2010 -87 2028 -62
rect 2073 -87 2091 -62
rect 2813 -45 2833 -15
rect 2864 -45 2884 -15
rect 3260 -87 3278 -62
rect 3323 -87 3341 -62
<< pdiffc >>
rect -823 248 -805 273
rect -731 160 -713 185
rect -418 248 -400 273
rect -326 160 -308 185
rect -6 136 14 166
rect 45 136 65 166
rect 332 248 350 273
rect 424 160 442 185
rect 680 248 698 273
rect 772 160 790 185
rect 1164 147 1184 177
rect 1215 147 1235 177
rect 1643 136 1663 166
rect 1694 136 1714 166
rect 1981 248 1999 273
rect 2073 160 2091 185
rect 2329 248 2347 273
rect 2421 160 2439 185
rect 2813 157 2833 187
rect 2864 157 2884 187
rect 3231 248 3249 273
rect 3323 160 3341 185
<< psubdiff >>
rect -65 41 -10 61
rect -65 11 -50 41
rect -30 11 -10 41
rect -65 1 -10 11
rect -842 -62 -802 -55
rect -842 -87 -829 -62
rect -811 -87 -802 -62
rect -842 -97 -802 -87
rect -437 -62 -397 -55
rect -437 -87 -424 -62
rect -406 -87 -397 -62
rect -437 -97 -397 -87
rect 661 -10 701 -3
rect 661 -35 674 -10
rect 692 -35 701 -10
rect 661 -45 701 -35
rect 1084 -13 1160 5
rect 1104 -43 1160 -13
rect 313 -62 353 -55
rect 313 -87 326 -62
rect 344 -87 353 -62
rect 313 -97 353 -87
rect 1084 -55 1160 -43
rect 1584 -22 1639 -2
rect 1584 -52 1599 -22
rect 1619 -52 1639 -22
rect 1584 -62 1639 -52
rect 2310 -10 2350 -3
rect 2310 -35 2323 -10
rect 2341 -35 2350 -10
rect 2310 -45 2350 -35
rect 2733 -13 2809 5
rect 2753 -43 2809 -13
rect 1962 -62 2002 -55
rect 1962 -87 1975 -62
rect 1993 -87 2002 -62
rect 1962 -97 2002 -87
rect 2733 -55 2809 -43
rect 3212 -62 3252 -55
rect 3212 -87 3225 -62
rect 3243 -87 3252 -62
rect 3212 -97 3252 -87
<< nsubdiff >>
rect -873 273 -832 285
rect -873 248 -861 273
rect -843 248 -832 273
rect -873 150 -832 248
rect -468 273 -427 285
rect -468 248 -456 273
rect -438 248 -427 273
rect -468 150 -427 248
rect -65 166 -10 306
rect -65 136 -50 166
rect -30 136 -10 166
rect -65 126 -10 136
rect 282 273 323 285
rect 282 248 294 273
rect 312 248 323 273
rect 282 150 323 248
rect 630 273 671 285
rect 630 248 642 273
rect 660 248 671 273
rect 630 150 671 248
rect 1079 255 1160 317
rect 1079 225 1088 255
rect 1108 225 1160 255
rect 1079 137 1160 225
rect 1584 166 1639 306
rect 1584 136 1599 166
rect 1619 136 1639 166
rect 1584 126 1639 136
rect 1931 273 1972 285
rect 1931 248 1943 273
rect 1961 248 1972 273
rect 1931 150 1972 248
rect 2279 273 2320 285
rect 2279 248 2291 273
rect 2309 248 2320 273
rect 2279 150 2320 248
rect 2728 265 2809 327
rect 2728 235 2737 265
rect 2757 235 2809 265
rect 2728 147 2809 235
rect 3181 273 3222 285
rect 3181 248 3193 273
rect 3211 248 3222 273
rect 3181 150 3222 248
<< psubdiffcont >>
rect -50 11 -30 41
rect -829 -87 -811 -62
rect -424 -87 -406 -62
rect 674 -35 692 -10
rect 1084 -43 1104 -13
rect 326 -87 344 -62
rect 1599 -52 1619 -22
rect 2323 -35 2341 -10
rect 2733 -43 2753 -13
rect 1975 -87 1993 -62
rect 3225 -87 3243 -62
<< nsubdiffcont >>
rect -861 248 -843 273
rect -456 248 -438 273
rect -50 136 -30 166
rect 294 248 312 273
rect 642 248 660 273
rect 1088 225 1108 255
rect 1599 136 1619 166
rect 1943 248 1961 273
rect 2291 248 2309 273
rect 2737 235 2757 265
rect 3193 248 3211 273
<< poly >>
rect 6 350 52 361
rect 6 332 17 350
rect 39 332 52 350
rect 6 324 52 332
rect 1190 351 1388 366
rect -759 285 -744 309
rect -354 285 -339 309
rect 20 306 35 324
rect 1190 317 1205 351
rect 1357 341 1406 351
rect -849 45 -804 59
rect -759 45 -744 150
rect -849 20 -842 45
rect -817 27 -744 45
rect -817 20 -804 27
rect -849 12 -804 20
rect -759 -55 -744 27
rect -444 45 -399 59
rect -354 45 -339 150
rect 396 285 411 309
rect 744 285 759 309
rect 20 111 35 126
rect 20 61 35 74
rect -444 20 -437 45
rect -412 27 -339 45
rect -412 20 -399 27
rect -444 12 -399 20
rect -354 -55 -339 27
rect 306 45 351 59
rect 396 45 411 150
rect 306 20 313 45
rect 338 27 411 45
rect 338 20 351 27
rect 306 12 351 20
rect 20 -28 35 1
rect 10 -35 45 -28
rect 10 -53 18 -35
rect 37 -53 45 -35
rect 10 -58 45 -53
rect 396 -55 411 27
rect 744 77 759 150
rect 1357 314 1367 341
rect 1395 314 1406 341
rect 2839 345 3005 360
rect 1357 303 1406 314
rect 1669 331 1848 339
rect 1669 324 1823 331
rect 1669 306 1684 324
rect 1815 314 1823 324
rect 1841 314 1848 331
rect 2839 327 2854 345
rect 2965 335 3005 345
rect 1190 122 1205 137
rect 1815 305 1848 314
rect 2045 285 2060 309
rect 2393 285 2408 309
rect 1669 111 1684 126
rect 781 89 823 97
rect 781 77 790 89
rect 744 67 790 77
rect 814 67 823 89
rect 744 62 823 67
rect 744 -3 759 62
rect 1955 45 2000 59
rect 2045 45 2060 150
rect 1955 20 1962 45
rect 1987 27 2060 45
rect 1987 20 2000 27
rect 1190 5 1205 18
rect 1955 12 2000 20
rect 744 -70 759 -45
rect 1669 -2 1684 11
rect 1326 -36 1373 -24
rect 1190 -66 1205 -55
rect 1326 -57 1337 -36
rect 1362 -57 1373 -36
rect 1326 -66 1373 -57
rect 2045 -55 2060 27
rect 2393 77 2408 150
rect 2965 317 2975 335
rect 2996 317 3005 335
rect 2965 312 3005 317
rect 3295 285 3310 309
rect 2839 132 2854 147
rect 2430 89 2472 97
rect 2430 77 2439 89
rect 2393 67 2439 77
rect 2463 67 2472 89
rect 2393 62 2472 67
rect 2393 -3 2408 62
rect 3205 45 3250 59
rect 3295 45 3310 150
rect 3205 20 3212 45
rect 3237 27 3310 45
rect 3237 20 3250 27
rect 2839 5 2854 18
rect 1190 -81 1373 -66
rect 1669 -83 1684 -62
rect 1736 -73 1776 -65
rect 1736 -83 1742 -73
rect 1669 -94 1742 -83
rect 1766 -94 1776 -73
rect -759 -122 -744 -97
rect -354 -122 -339 -97
rect 396 -122 411 -97
rect 1669 -98 1776 -94
rect 2393 -70 2408 -45
rect 2942 3 3004 20
rect 3205 12 3250 20
rect 2942 -21 2961 3
rect 2989 -21 3004 3
rect 2942 -37 3004 -21
rect 2839 -64 2854 -55
rect 2942 -64 2959 -37
rect 3295 -55 3310 27
rect 2839 -79 2959 -64
rect 1736 -103 1776 -98
rect 2045 -122 2060 -97
rect 3295 -118 3310 -97
<< polycont >>
rect 17 332 39 350
rect -842 20 -817 45
rect -437 20 -412 45
rect 313 20 338 45
rect 18 -53 37 -35
rect 1367 314 1395 341
rect 1823 314 1841 331
rect 790 67 814 89
rect 1962 20 1987 45
rect 1337 -57 1362 -36
rect 2975 317 2996 335
rect 2439 67 2463 89
rect 3212 20 3237 45
rect 1742 -94 1766 -73
rect 2961 -21 2989 3
<< locali >>
rect -849 285 -830 383
rect -445 285 -421 383
rect -55 306 -38 385
rect 6 350 52 361
rect 6 332 17 350
rect 39 332 52 350
rect 6 324 52 332
rect -872 273 -798 285
rect -872 248 -861 273
rect -843 248 -823 273
rect -805 248 -798 273
rect -872 240 -798 248
rect -467 273 -393 285
rect -467 248 -456 273
rect -438 248 -418 273
rect -400 248 -393 273
rect -467 240 -393 248
rect -739 185 -704 190
rect -739 160 -731 185
rect -713 160 -704 185
rect -739 150 -704 160
rect -334 185 -299 190
rect -334 160 -326 185
rect -308 160 -299 185
rect -334 150 -299 160
rect -65 166 -30 306
rect -848 45 -806 59
rect -848 20 -842 45
rect -817 20 -806 45
rect -848 12 -806 20
rect -730 44 -712 150
rect -324 149 -302 150
rect -443 45 -401 59
rect -730 40 -604 44
rect -730 23 -641 40
rect -617 23 -604 40
rect -730 19 -604 23
rect -443 20 -437 45
rect -412 20 -401 45
rect -730 -55 -712 19
rect -443 12 -401 20
rect -324 39 -306 149
rect -65 136 -50 166
rect -65 126 -30 136
rect -6 166 15 306
rect 14 136 15 166
rect -6 126 15 136
rect 39 166 70 306
rect 308 285 329 382
rect 662 285 682 384
rect 283 273 357 285
rect 283 248 294 273
rect 312 248 332 273
rect 350 248 357 273
rect 283 240 357 248
rect 631 273 705 285
rect 631 248 642 273
rect 660 248 680 273
rect 698 248 705 273
rect 631 240 705 248
rect 1085 255 1110 383
rect 1594 382 1612 385
rect 1357 342 1406 351
rect 1357 313 1365 342
rect 1397 313 1406 342
rect 1357 303 1406 313
rect 1594 306 1611 382
rect 1815 332 1848 339
rect 1815 313 1823 332
rect 1842 313 1848 332
rect 39 136 45 166
rect 65 136 70 166
rect 39 126 70 136
rect 375 214 565 231
rect -3 102 14 126
rect -152 85 14 102
rect -152 39 -133 85
rect -3 61 14 85
rect 45 102 62 126
rect 375 102 392 214
rect 416 185 451 190
rect 416 160 424 185
rect 442 160 451 185
rect 416 150 451 160
rect 45 85 392 102
rect 45 61 62 85
rect -324 21 -133 39
rect -65 41 -30 61
rect -324 -55 -306 21
rect -65 11 -50 41
rect -65 1 -30 11
rect -6 41 15 61
rect 14 11 15 41
rect -6 1 15 11
rect 39 41 70 61
rect 319 59 336 85
rect 39 11 45 41
rect 65 11 70 41
rect 307 45 349 59
rect 307 20 313 45
rect 338 20 349 45
rect 307 12 349 20
rect 425 39 448 150
rect 545 136 565 214
rect 725 220 986 237
rect 725 136 742 220
rect 764 185 799 190
rect 764 160 772 185
rect 790 170 799 185
rect 790 160 901 170
rect 764 150 901 160
rect 545 118 742 136
rect 781 89 823 97
rect 781 87 790 89
rect 694 67 790 87
rect 814 67 823 89
rect 694 66 823 67
rect 694 40 715 66
rect 781 62 823 66
rect 880 73 901 150
rect 968 119 986 220
rect 1085 225 1088 255
rect 1108 225 1110 255
rect 1169 253 1289 254
rect 1085 137 1110 225
rect 1128 236 1289 253
rect 1128 119 1145 236
rect 1164 177 1185 186
rect 1184 147 1185 177
rect 1164 137 1185 147
rect 1209 177 1240 186
rect 1209 147 1215 177
rect 1235 147 1240 177
rect 1209 137 1240 147
rect 968 102 1145 119
rect 1167 73 1184 137
rect 880 56 1184 73
rect 694 39 780 40
rect 425 21 780 39
rect 39 1 70 11
rect -842 -62 -767 -55
rect -842 -87 -829 -62
rect -811 -87 -794 -62
rect -776 -87 -767 -62
rect -842 -97 -767 -87
rect -739 -62 -704 -55
rect -739 -87 -731 -62
rect -713 -87 -704 -62
rect -739 -97 -704 -87
rect -437 -62 -362 -55
rect -437 -87 -424 -62
rect -406 -87 -389 -62
rect -371 -87 -362 -62
rect -437 -97 -362 -87
rect -334 -62 -299 -55
rect -334 -87 -326 -62
rect -308 -87 -299 -62
rect -334 -97 -299 -87
rect -815 -136 -792 -97
rect -407 -136 -389 -97
rect -55 -136 -38 1
rect 10 -35 45 -16
rect 425 -21 448 21
rect 10 -53 18 -35
rect 37 -53 45 -35
rect 10 -58 45 -53
rect 424 -55 448 -21
rect 661 -10 736 -3
rect 661 -35 674 -10
rect 692 -35 709 -10
rect 727 -35 736 -10
rect 661 -45 736 -35
rect 313 -62 388 -55
rect 313 -87 326 -62
rect 344 -87 361 -62
rect 379 -87 388 -62
rect 313 -97 388 -87
rect 416 -62 451 -55
rect 416 -87 424 -62
rect 442 -87 451 -62
rect 416 -97 451 -87
rect 345 -137 362 -97
rect 691 -134 708 -45
rect 759 -73 780 21
rect 797 -10 832 -3
rect 797 -35 805 -10
rect 823 -15 832 -10
rect 880 -15 901 56
rect 960 36 1140 39
rect 823 -35 901 -15
rect 959 22 1140 36
rect 797 -45 832 -35
rect 959 -73 978 22
rect 1084 -13 1104 5
rect 1084 -55 1104 -43
rect 759 -91 978 -73
rect 1085 -135 1102 -55
rect 1121 -91 1140 22
rect 1167 5 1184 56
rect 1215 113 1232 137
rect 1272 113 1289 236
rect 1584 166 1619 306
rect 1584 136 1599 166
rect 1584 126 1619 136
rect 1643 166 1664 306
rect 1663 136 1664 166
rect 1643 126 1664 136
rect 1688 166 1719 306
rect 1815 305 1848 313
rect 1952 285 1978 383
rect 2308 285 2333 383
rect 1932 273 2006 285
rect 1932 248 1943 273
rect 1961 248 1981 273
rect 1999 248 2006 273
rect 1932 240 2006 248
rect 2280 273 2354 285
rect 2280 248 2291 273
rect 2309 248 2329 273
rect 2347 248 2354 273
rect 2280 240 2354 248
rect 2734 265 2759 385
rect 2965 335 3005 345
rect 2965 317 2975 335
rect 2996 317 3005 335
rect 2965 312 3005 317
rect 3202 285 3228 384
rect 2374 237 2591 238
rect 2194 234 2214 235
rect 1688 136 1694 166
rect 1714 136 1719 166
rect 1688 126 1719 136
rect 2024 214 2214 234
rect 2024 213 2063 214
rect 1215 96 1289 113
rect 1646 102 1663 126
rect 1215 5 1232 96
rect 1497 85 1663 102
rect 1497 41 1516 85
rect 1431 39 1516 41
rect 1429 21 1516 39
rect 1164 -15 1185 5
rect 1184 -45 1185 -15
rect 1164 -55 1185 -45
rect 1209 -15 1240 5
rect 1209 -45 1215 -15
rect 1235 -45 1240 -15
rect 1209 -55 1240 -45
rect 1326 -36 1373 -24
rect 1326 -57 1337 -36
rect 1362 -57 1373 -36
rect 1326 -66 1373 -57
rect 1430 -91 1451 21
rect 1646 -2 1663 85
rect 1694 102 1711 126
rect 2024 102 2044 213
rect 2065 185 2100 190
rect 2065 160 2073 185
rect 2091 160 2100 185
rect 2065 150 2100 160
rect 2073 117 2097 150
rect 2194 136 2214 214
rect 2374 220 2635 237
rect 2374 136 2394 220
rect 2591 218 2635 220
rect 2413 185 2448 190
rect 2413 160 2421 185
rect 2439 170 2448 185
rect 2439 160 2550 170
rect 2413 150 2550 160
rect 2194 118 2394 136
rect 1694 85 2044 102
rect 1694 -2 1711 85
rect 1966 60 1987 85
rect 1956 45 1998 60
rect 1956 20 1962 45
rect 1987 20 1998 45
rect 1956 12 1998 20
rect 2074 39 2097 117
rect 2430 89 2472 97
rect 2430 87 2439 89
rect 2343 67 2439 87
rect 2463 67 2472 89
rect 2343 66 2472 67
rect 2343 40 2364 66
rect 2430 62 2472 66
rect 2529 91 2550 150
rect 2617 129 2635 218
rect 2734 235 2737 265
rect 2757 235 2759 265
rect 3182 273 3256 285
rect 2818 263 2938 264
rect 2734 147 2759 235
rect 2777 246 2938 263
rect 2777 129 2794 246
rect 2813 187 2834 196
rect 2833 157 2834 187
rect 2813 147 2834 157
rect 2858 187 2889 196
rect 2858 157 2864 187
rect 2884 157 2889 187
rect 2858 147 2889 157
rect 2617 113 2794 129
rect 2618 112 2794 113
rect 2816 91 2833 147
rect 2529 66 2833 91
rect 2343 39 2429 40
rect 2074 21 2429 39
rect 1584 -22 1619 -2
rect 1584 -52 1599 -22
rect 1584 -62 1619 -52
rect 1643 -22 1664 -2
rect 1663 -52 1664 -22
rect 1643 -62 1664 -52
rect 1688 -22 1719 -2
rect 2074 -21 2097 21
rect 2343 19 2364 21
rect 1688 -52 1694 -22
rect 1714 -52 1719 -22
rect 1688 -62 1719 -52
rect 2073 -55 2097 -21
rect 2310 -10 2385 -3
rect 2310 -35 2323 -10
rect 2341 -35 2358 -10
rect 2376 -35 2385 -10
rect 2310 -45 2385 -35
rect 1962 -62 2037 -55
rect 1121 -108 1451 -91
rect 1069 -138 1106 -135
rect 1594 -137 1611 -62
rect 1736 -73 1776 -65
rect 1736 -94 1742 -73
rect 1766 -94 1776 -73
rect 1736 -103 1776 -94
rect 1962 -87 1975 -62
rect 1993 -87 2010 -62
rect 2028 -87 2037 -62
rect 1962 -97 2037 -87
rect 2065 -62 2100 -55
rect 2065 -87 2073 -62
rect 2091 -87 2100 -62
rect 2065 -97 2100 -87
rect 1992 -137 2010 -97
rect 2333 -135 2356 -45
rect 2408 -73 2429 21
rect 2446 -10 2481 -3
rect 2446 -35 2454 -10
rect 2472 -15 2481 -10
rect 2529 -15 2550 66
rect 2609 36 2789 39
rect 2472 -35 2550 -15
rect 2608 22 2789 36
rect 2446 -45 2481 -35
rect 2608 -73 2627 22
rect 2733 -13 2753 5
rect 2733 -55 2753 -43
rect 2408 -91 2627 -73
rect 2734 -135 2751 -55
rect 2770 -92 2789 22
rect 2816 5 2833 66
rect 2864 123 2881 147
rect 2921 123 2938 246
rect 3182 248 3193 273
rect 3211 248 3231 273
rect 3249 248 3256 273
rect 3182 240 3256 248
rect 3315 185 3350 190
rect 3315 160 3323 185
rect 3341 160 3350 185
rect 3315 150 3350 160
rect 2864 106 2938 123
rect 2864 5 2881 106
rect 3206 45 3248 59
rect 3206 41 3212 45
rect 3077 21 3212 41
rect 2813 -15 2834 5
rect 2833 -45 2834 -15
rect 2813 -55 2834 -45
rect 2858 -15 2889 5
rect 2858 -45 2864 -15
rect 2884 -45 2889 -15
rect 2942 3 3004 20
rect 2942 -22 2961 3
rect 2989 -22 3004 3
rect 2942 -37 3004 -22
rect 2858 -55 2889 -45
rect 3077 -92 3095 21
rect 3206 20 3212 21
rect 3237 20 3248 45
rect 3206 12 3248 20
rect 3324 39 3345 150
rect 3324 21 3426 39
rect 3324 -55 3345 21
rect 2770 -111 3095 -92
rect 3212 -62 3287 -55
rect 3212 -87 3225 -62
rect 3243 -87 3260 -62
rect 3278 -87 3287 -62
rect 3212 -97 3287 -87
rect 3315 -62 3350 -55
rect 3315 -87 3323 -62
rect 3341 -87 3350 -62
rect 3315 -97 3350 -87
rect 2330 -136 2365 -135
rect 1069 -162 1070 -138
rect 1105 -162 1106 -138
rect 2330 -162 2365 -160
rect 2718 -138 2753 -135
rect 3241 -138 3260 -97
<< viali >>
rect -857 383 -822 407
rect -452 383 -417 407
rect -70 385 -35 409
rect 299 382 334 406
rect 653 384 688 408
rect -641 23 -617 40
rect 1079 383 1114 407
rect 1583 385 1618 409
rect 1948 383 1983 407
rect 2299 383 2334 407
rect 2728 385 2763 409
rect 1365 341 1397 342
rect 1365 314 1367 341
rect 1367 314 1395 341
rect 1395 314 1397 341
rect 1365 313 1397 314
rect 1823 331 1842 332
rect 1823 314 1841 331
rect 1841 314 1842 331
rect 1823 313 1842 314
rect 18 -53 37 -35
rect -821 -160 -786 -136
rect -416 -160 -381 -136
rect -66 -160 -31 -136
rect 336 -161 371 -137
rect 677 -158 712 -134
rect 3195 384 3230 408
rect 2961 -21 2989 3
rect 2961 -22 2989 -21
rect 1070 -162 1105 -138
rect 1585 -161 1620 -137
rect 1983 -161 2016 -137
rect 2330 -160 2365 -136
rect 2718 -162 2753 -138
rect 3233 -162 3268 -138
<< metal1 >>
rect -942 409 3429 413
rect -942 407 -70 409
rect -942 383 -857 407
rect -822 383 -452 407
rect -417 385 -70 407
rect -35 408 1583 409
rect -35 406 653 408
rect -35 385 299 406
rect -417 383 299 385
rect -942 382 299 383
rect 334 384 653 406
rect 688 407 1583 408
rect 688 384 1079 407
rect 334 383 1079 384
rect 1114 385 1583 407
rect 1618 407 2728 409
rect 1618 385 1948 407
rect 1114 383 1948 385
rect 1983 383 2299 407
rect 2334 385 2728 407
rect 2763 408 3429 409
rect 2763 385 3195 408
rect 2334 384 3195 385
rect 3230 384 3429 408
rect 2334 383 3429 384
rect 334 382 3429 383
rect -942 378 3429 382
rect 1356 342 1406 351
rect 1356 313 1365 342
rect 1397 313 1406 342
rect 1356 303 1406 313
rect 1815 332 1848 339
rect 1815 313 1823 332
rect 1842 313 1848 332
rect 1815 305 1848 313
rect -650 40 -580 44
rect -650 23 -641 40
rect -617 23 -580 40
rect -650 19 -580 23
rect -604 -16 -580 19
rect 1372 -16 1392 303
rect 1822 -16 1841 305
rect 2942 3 3004 20
rect 2942 -16 2961 3
rect -604 -22 2961 -16
rect 2989 -22 3004 3
rect -604 -33 3004 -22
rect 10 -35 45 -33
rect 10 -53 18 -35
rect 37 -53 45 -35
rect 2942 -37 3004 -33
rect 10 -58 45 -53
rect -945 -134 3441 -131
rect -945 -136 677 -134
rect -945 -160 -821 -136
rect -786 -160 -416 -136
rect -381 -160 -66 -136
rect -31 -137 677 -136
rect -31 -160 336 -137
rect -945 -161 336 -160
rect 371 -158 677 -137
rect 712 -136 3441 -134
rect 712 -137 2330 -136
rect 712 -138 1585 -137
rect 712 -158 1070 -138
rect 371 -161 1070 -158
rect -945 -162 1070 -161
rect 1105 -161 1585 -138
rect 1620 -161 1983 -137
rect 2016 -160 2330 -137
rect 2365 -138 3441 -136
rect 2365 -160 2718 -138
rect 2016 -161 2718 -160
rect 1105 -162 2718 -161
rect 2753 -162 3233 -138
rect 3268 -162 3441 -138
rect -945 -165 3441 -162
<< labels >>
rlabel metal1 -608 385 -553 406 1 vdd
port 1 n
rlabel polycont -437 20 -412 44 1 input
port 2 n
rlabel locali 3386 24 3415 36 1 output
port 3 n
rlabel locali -842 22 -816 46 1 Clk_in
port 4 n
rlabel metal1 -606 -160 -557 -138 1 vss
port 5 n
rlabel polycont 17 332 39 350 1 Clk_in
port 4 n
rlabel locali 1338 -58 1362 -36 1 Clk_in
port 4 n
rlabel polycont 1743 -93 1766 -74 1 Clk_in
port 4 n
rlabel locali 2975 317 2998 336 1 Clk_in
port 4 n
<< end >>
