module buffer (
    input wire in,    // Single input
    output wire out   // Single output
);

    // Assign the input to the output
    assign out = in;

endmodule