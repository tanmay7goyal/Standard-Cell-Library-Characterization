VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO D_FlipFlop_PosEdge
  CLASS BLOCK ;
  FOREIGN D_FlipFlop_PosEdge ;
  ORIGIN 9.450 1.650 ;
  SIZE 43.860 BY 5.780 ;
  PIN vdd
    ANTENNADIFFAREA 15.669000 ;
    PORT
      LAYER nwell ;
        RECT 27.100 3.450 28.270 3.460 ;
        RECT -8.920 1.180 -6.780 3.120 ;
        RECT -4.870 1.180 -2.730 3.120 ;
        RECT -0.850 1.060 1.240 3.240 ;
        RECT 2.630 1.180 4.770 3.120 ;
        RECT 6.110 1.180 8.250 3.120 ;
        RECT 10.610 1.170 12.940 3.350 ;
        RECT 15.640 1.060 17.730 3.240 ;
        RECT 19.120 1.180 21.260 3.120 ;
        RECT 22.600 1.180 24.740 3.120 ;
        RECT 27.100 1.270 29.430 3.450 ;
        RECT 31.620 1.180 33.760 3.120 ;
      LAYER li1 ;
        RECT -8.570 3.830 -8.220 4.070 ;
        RECT -4.520 3.830 -4.170 4.070 ;
        RECT -0.700 3.850 -0.350 4.090 ;
        RECT -8.490 2.850 -8.300 3.830 ;
        RECT -4.450 2.850 -4.210 3.830 ;
        RECT -0.550 3.060 -0.380 3.850 ;
        RECT 2.990 3.820 3.340 4.060 ;
        RECT 6.530 3.840 6.880 4.080 ;
        RECT -8.720 2.400 -7.980 2.850 ;
        RECT -4.670 2.400 -3.930 2.850 ;
        RECT -0.650 1.260 -0.300 3.060 ;
        RECT 3.080 2.850 3.290 3.820 ;
        RECT 6.620 2.850 6.820 3.840 ;
        RECT 10.790 3.830 11.140 4.070 ;
        RECT 15.830 3.850 16.180 4.090 ;
        RECT 2.830 2.400 3.570 2.850 ;
        RECT 6.310 2.400 7.050 2.850 ;
        RECT 10.850 1.370 11.100 3.830 ;
        RECT 15.940 3.820 16.120 3.850 ;
        RECT 19.480 3.830 19.830 4.070 ;
        RECT 22.990 3.830 23.340 4.070 ;
        RECT 27.280 3.850 27.630 4.090 ;
        RECT 15.940 3.060 16.110 3.820 ;
        RECT 15.840 1.260 16.190 3.060 ;
        RECT 19.520 2.850 19.780 3.830 ;
        RECT 23.080 2.850 23.330 3.830 ;
        RECT 19.320 2.400 20.060 2.850 ;
        RECT 22.800 2.400 23.540 2.850 ;
        RECT 27.340 1.470 27.590 3.850 ;
        RECT 31.950 3.840 32.300 4.080 ;
        RECT 32.020 2.850 32.280 3.840 ;
        RECT 31.820 2.400 32.560 2.850 ;
      LAYER met1 ;
        RECT -9.420 3.780 34.290 4.130 ;
    END
  END vdd
  PIN input
    ANTENNAGATEAREA 0.265500 ;
    PORT
      LAYER li1 ;
        RECT -4.430 0.120 -4.010 0.590 ;
    END
  END input
  PIN output
    ANTENNADIFFAREA 0.708000 ;
    PORT
      LAYER li1 ;
        RECT 33.150 1.500 33.500 1.900 ;
        RECT 33.240 0.390 33.450 1.500 ;
        RECT 33.240 0.210 34.260 0.390 ;
        RECT 33.240 -0.550 33.450 0.210 ;
        RECT 33.150 -0.970 33.500 -0.550 ;
    END
  END output
  PIN Clk_in
    ANTENNAGATEAREA 0.265500 ;
    PORT
      LAYER li1 ;
        RECT -8.480 0.120 -8.060 0.590 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.060 3.240 0.520 3.610 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.260 -0.660 13.730 -0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.360 -1.030 17.760 -0.650 ;
    END
    PORT
      LAYER li1 ;
        RECT 29.650 3.120 30.050 3.450 ;
    END
  END Clk_in
  PIN vss
    ANTENNADIFFAREA 4.012200 ;
    PORT
      LAYER li1 ;
        RECT -0.650 0.010 -0.300 0.610 ;
        RECT -8.420 -0.970 -7.670 -0.550 ;
        RECT -4.370 -0.970 -3.620 -0.550 ;
        RECT -8.150 -1.360 -7.920 -0.970 ;
        RECT -4.070 -1.360 -3.890 -0.970 ;
        RECT -0.550 -1.360 -0.380 0.010 ;
        RECT 6.610 -0.450 7.360 -0.030 ;
        RECT 3.130 -0.970 3.880 -0.550 ;
        RECT -8.210 -1.600 -7.860 -1.360 ;
        RECT -4.160 -1.600 -3.810 -1.360 ;
        RECT -0.660 -1.600 -0.310 -1.360 ;
        RECT 3.450 -1.370 3.620 -0.970 ;
        RECT 6.910 -1.340 7.080 -0.450 ;
        RECT 10.840 -0.550 11.040 0.050 ;
        RECT 3.360 -1.610 3.710 -1.370 ;
        RECT 6.770 -1.580 7.120 -1.340 ;
        RECT 10.850 -1.350 11.020 -0.550 ;
        RECT 15.840 -0.620 16.190 -0.020 ;
        RECT 23.100 -0.450 23.850 -0.030 ;
        RECT 10.690 -1.620 11.060 -1.350 ;
        RECT 15.940 -1.370 16.110 -0.620 ;
        RECT 19.620 -0.970 20.370 -0.550 ;
        RECT 19.920 -1.370 20.100 -0.970 ;
        RECT 23.330 -1.350 23.560 -0.450 ;
        RECT 27.330 -0.550 27.530 0.050 ;
        RECT 27.340 -1.350 27.510 -0.550 ;
        RECT 32.120 -0.970 32.870 -0.550 ;
        RECT 15.850 -1.610 16.200 -1.370 ;
        RECT 19.830 -1.610 20.160 -1.370 ;
        RECT 23.300 -1.620 23.650 -1.350 ;
        RECT 27.180 -1.620 27.530 -1.350 ;
        RECT 32.410 -1.380 32.600 -0.970 ;
        RECT 32.330 -1.620 32.680 -1.380 ;
      LAYER met1 ;
        RECT -9.450 -1.650 34.410 -1.310 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT -7.390 1.500 -7.040 1.900 ;
        RECT -3.340 1.500 -2.990 1.900 ;
        RECT -7.300 0.440 -7.120 1.500 ;
        RECT -3.240 1.490 -3.020 1.500 ;
        RECT -7.300 0.190 -6.040 0.440 ;
        RECT -3.240 0.390 -3.060 1.490 ;
        RECT -0.060 1.260 0.150 3.060 ;
        RECT 0.390 1.260 0.700 3.060 ;
        RECT 13.570 3.030 14.060 3.510 ;
        RECT 11.690 2.530 12.890 2.540 ;
        RECT 3.750 2.140 5.650 2.310 ;
        RECT -0.030 1.020 0.140 1.260 ;
        RECT -1.520 0.850 0.140 1.020 ;
        RECT -1.520 0.390 -1.330 0.850 ;
        RECT -0.030 0.610 0.140 0.850 ;
        RECT 0.450 1.020 0.620 1.260 ;
        RECT 3.750 1.020 3.920 2.140 ;
        RECT 4.160 1.500 4.510 1.900 ;
        RECT 0.450 0.850 3.920 1.020 ;
        RECT 0.450 0.610 0.620 0.850 ;
        RECT -3.240 0.210 -1.330 0.390 ;
        RECT -7.300 -0.550 -7.120 0.190 ;
        RECT -3.240 -0.550 -3.060 0.210 ;
        RECT -0.060 0.010 0.150 0.610 ;
        RECT 0.390 0.010 0.700 0.610 ;
        RECT 3.190 0.590 3.360 0.850 ;
        RECT 3.070 0.120 3.490 0.590 ;
        RECT 4.250 0.390 4.480 1.500 ;
        RECT 5.450 1.360 5.650 2.140 ;
        RECT 7.250 2.200 9.860 2.370 ;
        RECT 7.250 1.360 7.420 2.200 ;
        RECT 7.640 1.700 7.990 1.900 ;
        RECT 7.640 1.500 9.010 1.700 ;
        RECT 5.450 1.180 7.420 1.360 ;
        RECT 7.810 0.870 8.230 0.970 ;
        RECT 6.940 0.660 8.230 0.870 ;
        RECT 6.940 0.400 7.150 0.660 ;
        RECT 7.810 0.620 8.230 0.660 ;
        RECT 8.800 0.730 9.010 1.500 ;
        RECT 9.680 1.190 9.860 2.200 ;
        RECT 11.280 2.360 12.890 2.530 ;
        RECT 11.280 1.190 11.450 2.360 ;
        RECT 11.640 1.370 11.850 1.860 ;
        RECT 12.090 1.370 12.400 1.860 ;
        RECT 9.680 1.020 11.450 1.190 ;
        RECT 11.670 0.730 11.840 1.370 ;
        RECT 8.800 0.560 11.840 0.730 ;
        RECT 6.940 0.390 7.800 0.400 ;
        RECT 4.250 0.210 7.800 0.390 ;
        RECT -7.390 -0.970 -7.040 -0.550 ;
        RECT -3.340 -0.970 -2.990 -0.550 ;
        RECT 0.100 -0.580 0.450 -0.160 ;
        RECT 4.250 -0.210 4.480 0.210 ;
        RECT 4.240 -0.550 4.480 -0.210 ;
        RECT 4.160 -0.970 4.510 -0.550 ;
        RECT 7.590 -0.730 7.800 0.210 ;
        RECT 7.970 -0.150 8.320 -0.030 ;
        RECT 8.800 -0.150 9.010 0.560 ;
        RECT 9.600 0.360 11.400 0.390 ;
        RECT 7.970 -0.350 9.010 -0.150 ;
        RECT 9.590 0.220 11.400 0.360 ;
        RECT 7.970 -0.450 8.320 -0.350 ;
        RECT 9.590 -0.730 9.780 0.220 ;
        RECT 7.590 -0.910 9.780 -0.730 ;
        RECT 11.210 -0.910 11.400 0.220 ;
        RECT 11.670 0.050 11.840 0.560 ;
        RECT 12.150 1.130 12.320 1.370 ;
        RECT 12.720 1.130 12.890 2.360 ;
        RECT 16.430 1.260 16.640 3.060 ;
        RECT 16.880 1.260 17.190 3.060 ;
        RECT 18.150 3.050 18.480 3.390 ;
        RECT 28.180 2.630 29.380 2.640 ;
        RECT 27.770 2.460 29.380 2.630 ;
        RECT 23.740 2.370 25.910 2.380 ;
        RECT 21.940 2.340 22.140 2.350 ;
        RECT 20.240 2.140 22.140 2.340 ;
        RECT 20.240 2.130 20.630 2.140 ;
        RECT 12.150 0.960 12.890 1.130 ;
        RECT 16.460 1.020 16.630 1.260 ;
        RECT 12.150 0.050 12.320 0.960 ;
        RECT 14.970 0.850 16.630 1.020 ;
        RECT 14.970 0.410 15.160 0.850 ;
        RECT 14.310 0.390 15.160 0.410 ;
        RECT 14.290 0.210 15.160 0.390 ;
        RECT 11.640 -0.550 11.850 0.050 ;
        RECT 12.090 -0.550 12.400 0.050 ;
        RECT 14.300 -0.910 14.510 0.210 ;
        RECT 16.460 -0.020 16.630 0.850 ;
        RECT 16.940 1.020 17.110 1.260 ;
        RECT 20.240 1.020 20.440 2.130 ;
        RECT 20.650 1.500 21.000 1.900 ;
        RECT 20.730 1.170 20.970 1.500 ;
        RECT 21.940 1.360 22.140 2.140 ;
        RECT 23.740 2.200 26.350 2.370 ;
        RECT 23.740 1.360 23.940 2.200 ;
        RECT 25.910 2.180 26.350 2.200 ;
        RECT 24.130 1.700 24.480 1.900 ;
        RECT 24.130 1.500 25.500 1.700 ;
        RECT 21.940 1.180 23.940 1.360 ;
        RECT 16.940 0.850 20.440 1.020 ;
        RECT 16.940 -0.020 17.110 0.850 ;
        RECT 19.660 0.600 19.870 0.850 ;
        RECT 19.560 0.120 19.980 0.600 ;
        RECT 20.740 0.390 20.970 1.170 ;
        RECT 24.300 0.870 24.720 0.970 ;
        RECT 23.430 0.660 24.720 0.870 ;
        RECT 23.430 0.400 23.640 0.660 ;
        RECT 24.300 0.620 24.720 0.660 ;
        RECT 25.290 0.910 25.500 1.500 ;
        RECT 26.170 1.290 26.350 2.180 ;
        RECT 27.770 1.290 27.940 2.460 ;
        RECT 28.130 1.470 28.340 1.960 ;
        RECT 28.580 1.470 28.890 1.960 ;
        RECT 26.170 1.130 27.940 1.290 ;
        RECT 26.180 1.120 27.940 1.130 ;
        RECT 28.160 0.910 28.330 1.470 ;
        RECT 25.290 0.660 28.330 0.910 ;
        RECT 23.430 0.390 24.290 0.400 ;
        RECT 20.740 0.210 24.290 0.390 ;
        RECT 16.430 -0.620 16.640 -0.020 ;
        RECT 16.880 -0.620 17.190 -0.020 ;
        RECT 20.740 -0.210 20.970 0.210 ;
        RECT 23.430 0.190 23.640 0.210 ;
        RECT 20.730 -0.550 20.970 -0.210 ;
        RECT 11.210 -1.080 14.510 -0.910 ;
        RECT 20.650 -0.970 21.000 -0.550 ;
        RECT 24.080 -0.730 24.290 0.210 ;
        RECT 24.460 -0.150 24.810 -0.030 ;
        RECT 25.290 -0.150 25.500 0.660 ;
        RECT 26.090 0.360 27.890 0.390 ;
        RECT 24.460 -0.350 25.500 -0.150 ;
        RECT 26.080 0.220 27.890 0.360 ;
        RECT 24.460 -0.450 24.810 -0.350 ;
        RECT 26.080 -0.730 26.270 0.220 ;
        RECT 24.080 -0.910 26.270 -0.730 ;
        RECT 27.700 -0.920 27.890 0.220 ;
        RECT 28.160 0.050 28.330 0.660 ;
        RECT 28.640 1.230 28.810 1.470 ;
        RECT 29.210 1.230 29.380 2.460 ;
        RECT 28.640 1.060 29.380 1.230 ;
        RECT 28.640 0.050 28.810 1.060 ;
        RECT 32.060 0.410 32.480 0.590 ;
        RECT 30.770 0.210 32.480 0.410 ;
        RECT 28.130 -0.550 28.340 0.050 ;
        RECT 28.580 -0.550 28.890 0.050 ;
        RECT 29.420 -0.370 30.040 0.200 ;
        RECT 30.770 -0.920 30.950 0.210 ;
        RECT 32.060 0.120 32.480 0.210 ;
        RECT 27.700 -1.110 30.950 -0.920 ;
      LAYER met1 ;
        RECT 13.560 3.030 14.060 3.510 ;
        RECT 18.150 3.050 18.480 3.390 ;
        RECT -6.500 0.190 -5.800 0.440 ;
        RECT -6.040 -0.160 -5.800 0.190 ;
        RECT 13.720 -0.160 13.920 3.030 ;
        RECT 18.220 -0.160 18.410 3.050 ;
        RECT 29.420 -0.160 30.040 0.200 ;
        RECT -6.040 -0.330 30.040 -0.160 ;
        RECT 0.100 -0.580 0.450 -0.330 ;
        RECT 29.420 -0.370 30.040 -0.330 ;
  END
END D_FlipFlop_PosEdge
END LIBRARY

