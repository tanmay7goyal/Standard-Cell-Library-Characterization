magic
tech sky130A
timestamp 1725446438
<< nwell >>
rect -138 774 48 958
rect 182 774 368 958
<< nmos >>
rect -25 660 -10 707
rect 295 660 310 707
<< pmos >>
rect -25 795 -10 935
rect 295 795 310 935
<< ndiff >>
rect -65 691 -25 707
rect -65 669 -57 691
rect -39 669 -25 691
rect -65 660 -25 669
rect -10 691 30 707
rect -10 669 4 691
rect 22 669 30 691
rect -10 660 30 669
rect 255 691 295 707
rect 255 669 263 691
rect 281 669 295 691
rect 255 660 295 669
rect 310 691 350 707
rect 310 669 324 691
rect 342 669 350 691
rect 310 660 350 669
<< pdiff >>
rect -65 831 -25 935
rect -65 809 -57 831
rect -39 809 -25 831
rect -65 795 -25 809
rect -10 831 30 935
rect -10 809 4 831
rect 22 809 30 831
rect -10 795 30 809
rect 255 831 295 935
rect 255 809 263 831
rect 281 809 295 831
rect 255 795 295 809
rect 310 831 350 935
rect 310 809 324 831
rect 342 809 350 831
rect 310 795 350 809
<< ndiffc >>
rect -57 669 -39 691
rect 4 669 22 691
rect 263 669 281 691
rect 324 669 342 691
<< pdiffc >>
rect -57 809 -39 831
rect 4 809 22 831
rect 263 809 281 831
rect 324 809 342 831
<< psubdiff >>
rect -120 691 -65 707
rect -120 669 -108 691
rect -90 669 -65 691
rect -120 660 -65 669
rect 200 691 255 707
rect 200 669 212 691
rect 230 669 255 691
rect 200 660 255 669
<< nsubdiff >>
rect -120 831 -65 935
rect -120 809 -108 831
rect -90 809 -65 831
rect -120 795 -65 809
rect 200 831 255 935
rect 200 809 212 831
rect 230 809 255 831
rect 200 795 255 809
<< psubdiffcont >>
rect -108 669 -90 691
rect 212 669 230 691
<< nsubdiffcont >>
rect -108 809 -90 831
rect 212 809 230 831
<< poly >>
rect -25 935 -10 955
rect 295 935 310 955
rect -240 766 -165 776
rect -240 725 -230 766
rect -180 757 -165 766
rect -25 757 -10 795
rect 295 776 310 795
rect -180 734 -10 757
rect -180 725 -165 734
rect -240 713 -165 725
rect -25 707 -10 734
rect 235 769 310 776
rect 235 740 244 769
rect 287 740 310 769
rect 235 731 310 740
rect 295 707 310 731
rect -25 641 -10 660
rect 295 640 310 660
<< polycont >>
rect -230 725 -180 766
rect 244 740 287 769
<< locali >>
rect -135 1048 51 1117
rect 154 1048 332 1117
rect -78 935 -46 1048
rect 241 935 273 1048
rect -120 831 -28 935
rect -120 809 -108 831
rect -90 809 -57 831
rect -39 809 -28 831
rect -120 795 -28 809
rect -7 831 30 935
rect -7 809 4 831
rect 22 809 30 831
rect -7 795 30 809
rect 200 831 292 935
rect 200 809 212 831
rect 230 809 263 831
rect 281 809 292 831
rect 200 795 292 809
rect 313 831 350 935
rect 313 809 324 831
rect 342 809 350 831
rect 313 795 350 809
rect 2 776 27 795
rect -260 766 -165 776
rect -260 725 -230 766
rect -180 725 -165 766
rect -260 713 -165 725
rect 2 769 295 776
rect 2 740 244 769
rect 287 740 295 769
rect 2 731 295 740
rect 322 755 341 795
rect 2 707 27 731
rect 322 730 449 755
rect 322 707 341 730
rect -120 691 -28 707
rect -120 669 -108 691
rect -90 669 -57 691
rect -39 669 -28 691
rect -120 660 -28 669
rect -7 691 30 707
rect -7 669 4 691
rect 22 669 30 691
rect -7 660 30 669
rect 200 691 292 707
rect 200 669 212 691
rect 230 669 263 691
rect 281 669 292 691
rect 200 660 292 669
rect 313 691 350 707
rect 313 669 324 691
rect 342 669 350 691
rect 313 660 350 669
rect -88 583 -56 660
rect 235 583 267 660
rect -157 547 47 583
rect -159 509 47 547
rect 151 509 344 583
<< viali >>
rect 51 1048 154 1117
rect 47 509 151 583
<< metal1 >>
rect -181 1117 372 1133
rect -181 1048 51 1117
rect 154 1048 372 1117
rect -181 1018 372 1048
rect -188 583 377 602
rect -188 509 47 583
rect 151 509 377 583
rect -188 487 377 509
<< labels >>
rlabel polycont -230 725 -183 764 1 in
port 1 n
rlabel locali 414 736 434 748 1 out2
port 2 n
rlabel metal1 227 1069 265 1098 1 vdd
port 3 n
rlabel metal1 200 532 238 561 1 gnd
port 4 n
<< end >>
